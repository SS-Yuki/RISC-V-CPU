// `ifndef __MUL_VALID_SV
// `define __MUL_VALID_SV

// `ifdef VERILATOR
// `include "include/common.sv"
// `include "include/pipes.sv"
// `else

// `endif


// module mul_valid
// 	import common::*;
// 	import pipes::*;(
// 	input u1 mulalu_type,
// 	input u1 finish,
// 	output u1 valid
// );
// 	assign valid = mulalu_
	
// endmodule

// `endif

